module adder(

input wire [31:0]IN1,
input wire [31:0]IN2,
output wire [31:0]OUT

);

assign OUT = IN1 + IN2 ;


endmodule







